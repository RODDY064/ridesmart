<?xml version="1.0" encoding="UTF-8"?>
<svg id="Layer_1" data-name="Layer 1" xmlns="http://www.w3.org/2000/svg" viewBox="0 0 450 450">
  <path d="M404.46,185.87c-1.24-7.38-2.91-13.92-5.17-17.72-.79-1.34-1.66-2.34-2.61-2.92h-.01c-.26-.16-.52-.29-.8-.37-.02,0-.03-.02-.05-.02-.05-.02-.1-.04-.15-.05H40.57s-9.21-3.07-7.67,44.51c.04,1.77,.07,3.47,.1,5.12,.35,19.33,.4,30.97,.33,37.99,0,1.06-.02,2.03-.04,2.89-.12,7.47-.39,7.74-.39,7.74,0,0,0,1.54,2.05,2.05,2.05,.51,4.69,0,4.69,0l21.41,3.58H127.92s-4.96-30.7,21.65-30.7c14.07,0,19.41,8.15,21.32,15.83,1.7,6.86,.68,13.33,.68,13.33l12.79,.14,131.49,1.4s-5.11-29.68,20.98-29.68,20.07,29.68,20.07,29.68h38.48s10.01-.69,12.57-4.18v-36.76s-.41-23.54-3.49-41.85h0ZM96.31,265.89v-4.27h9.6v4.27h-9.6Zm152.5,.2v-4.61h10.29v4.61h-10.29Z" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <polyline points="104.72 164.74 104.72 161.71 75.27 161.71 75.27 164.74" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <path d="M386.73,164.74v-2.31s4.1-.04,6.52,1.16c2.41,1.2,3.42,1.64,3.42,1.64" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <path d="M404.46,185.87h3.66c.83,0,1.55,.6,1.69,1.42,.5,2.84,1.5,9.4,1.15,14.85h6.7c.51-3.58,.83-9.8-2.05-16.37-.5-1.15-1.06-2.21-1.63-3.16-.54-.9-1.5-1.46-2.55-1.48l-7.84,.03" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <path d="M407.94,221.09h2.97s1.12,7.65-.93,12.26l-2.05,4.6" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <path d="M166.94,262s2-19.15-16.37-20.47c-21.49-1.53-19.83,20.47-19.83,20.47,0,0,.07,17.25,18.14,17.32,18.06,.08,18.06-17.32,18.06-17.32Z" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <polyline points="32.89 209.3 40.05 214.41 39.62 265.07" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <line x1="33.28" y1="255.29" x2="39.7" y2="255.29" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <line x1="32.89" y1="252.4" x2="40.05" y2="252.4" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <polyline points="33.28 217.55 43.56 217.56 184.34 218 184.34 235.05 43.63 234.88 43.63 218.51 42.61 218.51 42.61 234.37 41.59 234.37 41.59 218.51 40.05 218.44" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <polyline points="32.98 214.41 40.05 214.41 40.56 164.78" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <polygon points="43.63 238.46 43.63 263.31 50.75 263.31 50.75 265.07 58.58 265.07 58.58 265.89 82.54 265.89 82.54 238.46 43.63 238.46" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <polygon points="80.98 262 80.98 239.59 44.33 239.59 44.33 262.3 80.98 262" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <polygon points="117.27 238.46 117.27 265.89 105.92 265.89 105.92 261.62 96.31 261.62 96.31 265.89 83.91 265.89 83.91 238.46 117.27 238.46" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <polyline points="117.27 238.46 117.27 237.18 120.09 237.18 120.09 265.89 124.6 268.65" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <polyline points="184.34 267.25 184.34 237.58 146.99 236.42 170.87 237.27 170.87 253.8" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <path d="M149.04,251.77c.55,0,4.59,.19,7.16,3.58,2.47,3.25,1.66,6.95,1.54,7.68-1.02,6.14-5.63,9.21-10.74,8.7-5.84-.58-9.1-5.76-8.7-10.74,.24-2.99,1.62-7.17,5.12-8.7,2.37-1.06,4.62-.73,5.62-.52h0Z" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <path d="M149.04,257.39c2.44,.35,4.3,2.2,4.55,4.36,.33,2.87-2.3,5.23-4.73,5.5-1.55,.17-2.91-.26-3.91-1.1-1.3-1.08-2-2.81-1.77-4.4,.35-2.4,2.8-4.41,5.86-4.36Z" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <path d="M354.73,263.02s2-19.15-16.37-20.47c-21.49-1.54-19.83,20.47-19.83,20.47,0,0,.07,17.25,18.14,17.32,18.06,.08,18.06-17.32,18.06-17.32h0Z" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <path d="M336.82,252.79c.55,0,4.59,.19,7.16,3.58,2.47,3.25,1.69,6.95,1.54,7.67-.91,4.33-5.09,9.17-10.75,8.7-5.85-.49-9.51-6.35-9.11-11.33,.24-2.99,2.03-6.58,5.53-8.11,2.39-1.04,4.63-.72,5.63-.51h0Z" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <path d="M336.82,258.42c2.44,.35,4.3,2.2,4.55,4.36,.33,2.87-2.3,5.23-4.73,5.5-1.55,.17-2.91-.26-3.91-1.1-1.3-1.08-2-2.81-1.77-4.4,.35-2.41,2.8-4.42,5.86-4.36h0Z" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <polyline points="40.05 214.41 182.29 214.41 182.29 176.66 40.56 176.66" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <polyline points="40.46 174.86 391.7 174.65 391.7 164.74" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <polyline points="392.66 164.78 392.66 176.64 184.34 176.66 184.34 179.39 183.28 179.39 183.35 214.41 184.34 214.41 184.34 218" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <line x1="216.08" y1="176.66" x2="216.08" y2="214.41" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <polyline points="184.34 179.39 216.08 179.39 216.08 180.47 183.29 180.47" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <polygon points="215.11 214.41 214.02 216.46 214.02 218 347.19 218 362.4 223.11 362.4 219.32 352.17 215.44 360.87 215.44 360.89 214.41 215.11 214.41" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <polyline points="214.02 218 214.02 235.05 362.4 235.05 362.4 223.11" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <path d="M185.36,266.09v-48.54l-.09-3.14c-.6-.51-.93-1.73-.93-1.73v-28.45c0-2.55,2.5-2.56,2.5-2.56h25.13c1.03,0,1.54,1.09,1.54,1.09v29.61c0,1.02-1.23,2.05-1.23,2.05l.21,51.68h-27.13Z" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <rect x="187.25" y="185.99" width="23.89" height="28.43" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <polyline points="362.4 235.05 362.4 267.16 395.66 267.16 395.66 179.95 396.5 179.95 396.5 176.67 392.66 176.64" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <polyline points="361.89 219.02 361.89 180.69 395.66 180.69" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <line x1="360.87" y1="218.51" x2="360.87" y2="176.64" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <path d="M364.96,182.69h25.72s2.42,.51,2.93,3.07v79.82h-29.54v-78.82s-.65-3.05,.89-4.07Z" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <polygon points="390.03 227.72 390.03 187.58 366.64 187.58 366.64 221.9 390.03 227.72" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <path d="M366.64,224.14l20.69,5.33c1.59,.41,2.7,1.84,2.7,3.49v30.41l-21.33-.63c-1.15-.03-2.06-.98-2.06-2.13v-36.47h0Z" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <polyline points="63.06 176.66 63.06 214.41 64.56 214.41 64.61 188.32 116.8 188.32 116.8 214.41 118.68 214.41 118.68 176.66" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <rect x="66.66" y="181.67" width="48.19" height="5.5" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <rect x="234.48" y="178.6" width="43.28" height="7.65" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <polyline points="279.77 176.65 279.77 214.41 280.78 214.41 280.78 176.65" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <polyline points="311.49 176.65 311.49 214.41 312.5 214.41 312.5 176.65" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <path d="M399.29,168.15v54.23c-.05,4.31,1.59,6.4,4.28,8.3,1.16,.82,2.6,1.69,4.37,2.54" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <path d="M397.19,267.16s4.03-.02,6.84-1.79c1.49-.94,2.37-2.61,2.37-4.37v-17.79c0-2.22-1.03-4.31-2.77-5.68-2.03-1.6-5.93-2.14-6.44-2.48v32.11Z" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <rect x="96.31" y="261.62" width="9.6" height="4.27" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <polygon points="280.27 236.42 280.27 266.09 259.11 266.09 259.11 261.49 248.81 261.49 248.81 266.09 228.06 266.09 228.06 236.42 280.27 236.42" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <rect x="248.81" y="261.49" width="10.29" height="4.61" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <line x1="44.19" y1="261.09" x2="81.04" y2="261.09" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <line x1="44.19" y1="259.16" x2="81.04" y2="259.16" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <line x1="44.19" y1="257.22" x2="81.04" y2="257.22" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <line x1="44.19" y1="255.28" x2="81.04" y2="255.28" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <line x1="44.19" y1="253.34" x2="81.04" y2="253.34" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <line x1="44.19" y1="251.4" x2="81.04" y2="251.4" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <line x1="44.19" y1="249.46" x2="81.04" y2="249.46" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <line x1="44.19" y1="247.52" x2="81.04" y2="247.52" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <line x1="44.19" y1="245.58" x2="81.04" y2="245.58" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <line x1="44.19" y1="243.64" x2="81.04" y2="243.64" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
  <line x1="44.19" y1="241.7" x2="81.04" y2="241.7" fill="none" stroke="#000" stroke-miterlimit="10" stroke-width=".5"/>
</svg>